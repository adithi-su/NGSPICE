.include ./t14y_tsmc_025_level3.txt

*netlist
m0 out in 0 0 cmosn l=1.8u w=6.4u 
r0 vdd out 100

*power sources
Vdd vdd 0 5
Vin in 0 dc 2.5 pulse(0 5 0.01n 0.05n 0.05n 10n 20n) 

* computing the response for various load resistance values
.control
foreach res 100 1k 100k
alter r0=$res
tran 0.1ns 2n
dc Vin 0 5 0.1
end
.endc 

.control
foreach iter 1 2 3
setplot dc$iter
setplot tran$iter
end

plot tran1.in tran1.out tran2.out tran3.out
plot dc1.out dc2.out dc3.out vs in
plot tran1.Vdd#branch*vdd*-1 tran2.Vdd#branch*vdd*-1 tran3.Vdd#branch*vdd*-1
.endc
.end                                                                      
