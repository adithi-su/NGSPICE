* cmos inverter characteristics

* include the model files
.include ./t14y_tsmc_025_level3.txt
  
* netlist
* m_instance_name drain_node gate_node source_node bulk_substrate_node model_name L=length W=width
m1 out in 0 0 cmosn l=1u w=1u 
m2 out in vdd vdd cmosp l=1u w=2u


* power sources excitation etc.
* v_instance_name posive_node negetive_node value
v_dd vdd 0 3.3
v_in in 0 pulse(0 3.3 0 0.05n 0.05n 0.5n 1n)

.control
    tran 0.01n 2n
    setplot tran1
    plot in out
    plot -v_dd#branch
    dc v_in 0 3.3 0.1 
    setplot dc1
    plot in out
    plot -v_dd#branch
.endc

.end