.include ./t14y_tsmc_025_level3.txt
  
m1 out in 0 0 cmosn l=1u w=1u 
m2 out in vdd vdd cmosp l=1u w=2u

v_dd vdd 0 dc 5
v_in in 0 dc 5

.dc v_in 0 5 0.1

.control
run
plot out,in
.endc
.end
