* rc simulation

*rc time constant = 1ms
r0 in out 1
c0 out 0 1m

* pulse on period = 1e06 times rc time constant
Vin in 0 dc 2.5 pulse(0 1 1n 0.0001n 0.0001n 1 2) 

.op

.control
tran 0.1ms 10ms
setplot tran1
plot -vin#branch
plot in out in-out
.endc

.end
