.include ./t14y_tsmc_025_level3.txt

* F = (A.B)'  NAND

m1 F A int 0 cmosn L=1u W=10u
m2 int B 0 0 cmosn L=1u W=10u

m3 F A vdd vdd cmosp L=1u W=10u
m4 F B vdd vdd cmosp L=1u W=10u

v_dd vdd 0 3.3
v_1 A 0 PULSE(0 3.3 0 0 0 8ns 16ns)
v_2 B 0 PULSE(0 3.3 0 0 0 16ns 32ns)

.control
tran 0.1ns 32ns
run
end
plot tran1.A tran1.B tran1.F
.endc
.end
