.include ./t14y_tsmc_025_level3.txt

*netlist
m1 vdd in s 0 cmosn l=1u w=0.55u

*power sources
v_dd vdd 0 5
v_in in 0 5
v_ss s 0 0

.dc v_in 0 5 0.1 v_ss 0 3 1
.control
run
setplot dc1
plot -v_dd#branch
.endc
.end
				
